example-1.C MAXIMUM POWER TRANSFER THEOREM
V1 1 0 5
R1 1 2 2.2K
R2 2 4 1.2K
R3 1 3 4.7K
R4 3 0 3.5K
R5 3 4 2K
R6 4 0 3K
R7 4 5 2.5K
R8 5 0 {RLOAD}
.PARAM RLOAD=2K
.STEP PARAM RLOAD 1K 5K 100
.op

.END
