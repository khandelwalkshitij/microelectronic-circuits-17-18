EXAMPLE-5B SERIES RESONANCE
VIN 1 0 AC PULSE(0 5 0 10P 10P 0.5M 1M)
R1  1 2 10K
L1  2 3 1U
C1  3 0 0.01U
*.TRAN 0.1M 5M 0
.AC DEC 10 10MEG 10
.END
