EXAMPLE-7 NMOS MOSFET IV CHARACTERISTICS

*** 1.2um techbology level=3 MODEL file ****
.MODEL CMOSN  NMOS LEVEL=3 PHI=0.600000 TOX=2.1200E-08 XJ=0.200000U
+TPG=1 VTO=0.7860 DELTA=6.9670E-01 LD=1.6470E-07 KP=9.6379E-05
+UO=591.7 THETA=8.1220E-02 RSH=8.5450E+01 GAMMA=0.5863
+NSUB=2.7470E+16 NFS=1.98E+12 VMAX=1.7330E+05 ETA=4.3680E-02
+KAPPA=1.3960E-01 CGDO=4.0241E-10 CGSO=4.0241E-10
+CGBO=3.6144E-10 CJ=3.8541E-04 MJ=1.1854 CJSW=1.3940E-10
+MJSW=0.125195 PB=0.800000

M1 1 2 0 4 CMOSN L=1.2U W=6U
VGS 2 0 2.5
VDS 1 0 4.0
VBS 4 0 0

*.DC VDS 0 5 0.1 VGS 0 5 1 ; DC CAHRACTERISTICS
.DC VGS 0 5 0.1 VBS 0 -3 1 ; STUDY BODY EFFECT

.END
