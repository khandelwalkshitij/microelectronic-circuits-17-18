Example-2 PN Junction IV Characteristics
.MODEL PN1N4007 d(IS=7.02767e-09 RS=0.0341512 N=1.80803 EG=1.05743
+XTI=5 BV=1000 IBV=5e-08 CJO=1e-11
+VJ=0.7 M=0.5 FC=0.5 TT=1e-07
+KF=0 AF=1)

VA 1 0 5V
R1 1 2 470
D1 2 0 PN1N4007
*.DC VA 0 1.5 0.1 ;FORWARD BIAS CHARCTERISTICS
.DC VA 0 -2 0.01 TEMP 20 40 10 ;REVERSE BIAS CHARCTERISTICS WITH TEMPERATURE DEPENDENCE
.OP ; OPERATING POINT
.END
