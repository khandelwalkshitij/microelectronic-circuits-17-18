Example-4 PN Junction diode Clipper 
.MODEL DI_1N4007 D  ( IS=76.9p RS=42.0m BV=1.00k IBV=5.00u
+ CJO=26.5p  M=0.333 N=1.45 TT=4.32u )
VIN 1 0 SIN (0V 5V 1.0K)
R1 1 2 470
D1 2 3 DI_1N4007
VA 3 0 1.5V
D2 4 2 DI_1N4007
VB 4 0 -1.5V
.TRAN 0.01M 5M 0M
.END
