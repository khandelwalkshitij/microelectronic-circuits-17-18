Example-3 Zener diode VOLTAGE REGULATOR Chartacteristics

.SUBCKT BZX84C6V2_CS  1 2
*        Terminals    A   K
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 5.12
.MODEL DF D ( IS=23.3p RS=33.4 N=1.10
+ CJO=63.9p VJ=0.750 M=0.330 TT=50.1n )
.MODEL DR D ( IS=4.65f RS=2.30 N=1.49 )
.ENDS

VA 1 0 8

R1 1 2 100

X1 3 2 BZX84C6V2_CS ;ZENER DIODE

RL 2 0 {RLOAD}

VZ 3 0 0 ; ACTS LIKE AMMETER

.OP

*.DC VA 0 10 0.01 ; TO OBSERVE IV CHARCTERISTICS
.PARAM RLOAD=200
.STEP PARAM RLOAD 200 500 20
.END
