EXAMPLE-6 CE CONFIGURATION IV CAHRACTERISTICS BC107 
* ADDING MODEL FILE FOR BJT
*
.lib D:\myLib.lib
*
*------------NETLIST BEGINS HERE ---------------------*
VCC 1 0 5
VBB 3 0 5
Q1 1 2 0 BC107A
RB 3 2   100K

*----------------------- ANALYSIS BEGINS HERE ----------------*
.OP
.DC VCC 0 5 0.1 VBB 2 5 1 
.END