EXAMPLE-5B BAND PASS FILTER
VIN 1 0 AC sin(0 5 1k)
R1  1 2 200
C1  2 0 0.25u
C2  2 3 1U
R2  3 0 1.0K
.AC DEC 10 5k 100
.END
