EXAMPLE-6 CE CONFIGURATION IV CAHRACTERISTICS BC107 
* ADDING MODEL FILE FOR BJT
*
.model BC107A   NPN(Is=7.049f Xti=3 Eg=1.11 Vaf=116.3 Bf=375.5 Ise=7.049f
+               Ne=1.281 Ikf=4.589 Nk=.5 Xtb=1.5 Br=2.611 Isc=121.7p Nc=1.865
+               Ikr=5.313 Rc=1.464 Cjc=5.38p Mjc=.329 Vjc=.6218 Fc=.5 Cje=11.5p
+               Mje=.2717 Vje=.5 Tr=10n Tf=451p Itf=6.194 Xtf=17.43 Vtf=10)
*
*------------NETLIST BEGINS HERE ---------------------*
VCC 1 0 5
VBB 3 0 5
Q1 1 2 0 BC107A
RB 3 2   100K

*----------------------- ANALYSIS BEGINS HERE ----------------*
.OP
.DC VCC 0 5 0.1 VBB 2 5 1 
.END
